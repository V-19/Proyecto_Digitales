// 10'b1010010110; //D5.6 impar = 1010010110
// 10'b1001000101; 	//D16.2 impar = 1001000101
// 10'b1100000101;	// K28.5 par = 1100000101
// 10'b0011111010; //K28.5 impar = 0011111010
// 10'b1101101000; //K27.7 impar = 1101101000
// 10'b0010010111; //K27.7 par = 0010010111
// 10'b1001110100; //D0.0 impar = 1001110100\
// 10'b0110001011; //D0.0 par = 0110001011
// 10'b0111010100; //D1.0 impar = 0111010100
// 10'b1000101011;//D1.0 par = 1000101011
// 10'b1011010100;//D2.0 impar = 1011010100
// 10'b0100101011;//D2.0 par = 0100101011
// 10'b1100011011;//D3.0 impar = 1100011011
// 10'b1100010100;//D3.0 par = 1100010100
// 10'b1101010100;//D4.0 impar = 1101010100
// 10'b0010101011;//D4.0 par = 0010101011
// 10'b1010011011;//D5.0 impar = 1010011011
// 10'b1010010100;//D5.0 par = 1010010100
// 10'b0110011011;//D6.0 impar = 0110011011
// 10'b0110010100;//D6.0 par = 0110010100
// 10'b1110001011;//D7.0 impar = 1110001011
// 10'b0001110100;//D7.0 par = 0001110100
// 10'b0001101011;//D8.0 par = 0001101011
// 10'b1110010100;//D8.0 impar = 1110010100
// 10'b1001011011;//D9.0 impar = 1001011011
// 10'b1001010100;//D9.0 par = 1001010100
// 10'b0100010111;//K29.7 = 0100010111 par
// 10'b1011101000;//K29.7 = 1011101000 impar

//hex		//binary
//I/ IDLE 1 //K28.5/D5.6
//I/ IDLE 2 //K28.5/D16.2
module cgroup(tx_octect,
              code_group_Imp,
              code_group_Par,
              );
    
    output reg [7:0]tx_octect[267:0]     ; //8'b10101111;//R/K23.7
    output reg [9:0]code_group_Imp[267:0];  //8'b11111011; //S/k27.7
    output reg [9:0]code_group_Par[267:0];  //8'b11111101;  //T/K29.7
                                            // reg [9:0] code_group [0:27][1:0];
    
    
    // code_group[0][0] = 10'b0000000001;
    // code_group[0][1] = 10'b1010010110;  //D5.6 impar = 1010010110
    // code_group[1][0] = 10'b1001000101; 	//D16.2 impar = 1001000101
    // code_group[2][0] = 10'b1100000101;	 // K28.5 par = 1100000101
    // code_group[3][0]  = 10'b0011111010;  //K28.5 impar  = 0011111010
    // code_group[4][0]  = 10'b1101101000;  //K27.7 impar  = 1101101000
    // code_group[5][0]  = 10'b0010010111;  //K27.7 par  = 0010010111
    // code_group[6][0]  = 10'b1001110100;  //D0.0 impar  = 1001110100\
    // code_group[7][0]  = 10'b0110001011;  //D0.0 par  = 0110001011
    // code_group[8][0]  = 10'b0111010100;  //D1.0 impar  = 0111010100
    // code_group[9][0]  = 10'b1000101011;  //D1.0 par  = 1000101011
    // code_group[10][0] = 10'b1011010100;  //D2.0 impar = 1011010100
    // code_group[11][0] = 10'b0100101011;  //D2.0 par = 0100101011
    // code_group[12][0] = 10'b1100011011;  //D3.0 impar = 1100011011
    // code_group[13][0] = 10'b1100010100;  //D3.0 par = 1100010100
    // code_group[14][0] = 10'b1101010100;  //D4.0 impar = 1101010100
    // code_group[15][0] = 10'b0010101011;  //D4.0 par = 0010101011
    // code_group[16][0] = 10'b1010011011;  //D5.0 impar = 1010011011
    // code_group[17][0] = 10'b1010010100;  //D5.0 par = 1010010100
    // code_group[18][0] = 10'b0110011011;  //D6.0 impar = 0110011011
    // code_group[19][0] = 10'b0110010100;  //D6.0 par = 0110010100
    // code_group[20][0] = 10'b1110001011;  //D7.0 impar = 1110001011
    // code_group[21][0] = 10'b0001110100;  //D7.0 par = 0001110100
    // code_group[22][0] = 10'b0001101011;  //D8.0 par = 0001101011
    // code_group[23][0] = 10'b1110010100;  //D8.0 impar = 1110010100
    // code_group[24][0] = 10'b1001011011;  //D9.0 impar = 1001011011
    // code_group[25][0] = 10'b1001010100;  //D9.0 par = 1001010100
    // code_group[26][0] = 10'b0100010111;  //K29.7 = 0100010111 par
    // code_group[27][0] = 10'b1011101000;  //K29.7 = 1011101000 impar
    
                                // assign code_r ;                                                                                                                                                                                          //R/K23.7
                                // assign code_s ;                                                                                                                                                                                          //S/k27.7
                                // assign code_t ;                                                                                                                                                                                          //T/K29.7
                                //V/30.7
    //Octect Values
    always begin
	tx_octect[0]   = 00000000; //Value before code_group
    tx_octect[1]   = 00000001; //Value before code_group
    tx_octect[2]   = 00000010; //Value before code_group
    tx_octect[3]   = 00000011; //Value before code_group
    tx_octect[4]   = 00000100; //Value before code_group
    tx_octect[5]   = 00000101; //Value before code_group
    tx_octect[6]   = 00000110; //Value before code_group
    tx_octect[7]   = 00000111; //Value before code_group
    tx_octect[8]   = 00001000; //Value before code_group
    tx_octect[9]   = 00001001; //Value before code_group
    tx_octect[10]  = 00001010; //Value before code_group
    tx_octect[11]  = 00001011; //Value before code_group
    tx_octect[12]  = 00001100; //Value before code_group
    tx_octect[13]  = 00001101; //Value before code_group
    tx_octect[14]  = 00001110; //Value before code_group
    tx_octect[15]  = 00001111; //Value before code_group
    tx_octect[16]  = 00010000; //Value before code_group
    tx_octect[17]  = 00010001; //Value before code_group
    tx_octect[18]  = 00010010; //Value before code_group
    tx_octect[19]  = 00010011; //Value before code_group
    tx_octect[20]  = 00010100; //Value before code_group
    tx_octect[21]  = 00010101; //Value before code_group
    tx_octect[22]  = 00010110; //Value before code_group
    tx_octect[23]  = 00010111; //Value before code_group
    tx_octect[24]  = 00011000; //Value before code_group
    tx_octect[25]  = 00011001; //Value before code_group
    tx_octect[26]  = 00011010; //Value before code_group
    tx_octect[27]  = 00011011; //Value before code_group
    tx_octect[28]  = 00011100; //Value before code_group
    tx_octect[29]  = 00011101; //Value before code_group
    tx_octect[30]  = 00011110; //Value before code_group
    tx_octect[31]  = 00011111; //Value before code_group
    tx_octect[32]  = 00100000; //Value before code_group
    tx_octect[33]  = 00100001; //Value before code_group
    tx_octect[34]  = 00100010; //Value before code_group
    tx_octect[35]  = 00100011; //Value before code_group
    tx_octect[36]  = 00100100; //Value before code_group
    tx_octect[37]  = 00100101; //Value before code_group
    tx_octect[38]  = 00100110; //Value before code_group
    tx_octect[39]  = 00100111; //Value before code_group
    tx_octect[40]  = 00101000; //Value before code_group
    tx_octect[41]  = 00101001; //Value before code_group
    tx_octect[42]  = 00101010; //Value before code_group
    tx_octect[43]  = 00101011; //Value before code_group
    tx_octect[44]  = 00101100; //Value before code_group
    tx_octect[45]  = 00101101; //Value before code_group
    tx_octect[46]  = 00101110; //Value before code_group
    tx_octect[47]  = 00101111; //Value before code_group
    tx_octect[48]  = 00110000; //Value before code_group
    tx_octect[49]  = 00110001; //Value before code_group
    tx_octect[50]  = 00110010; //Value before code_group
    tx_octect[51]  = 00110011; //Value before code_group
    tx_octect[52]  = 00110100; //Value before code_group
    tx_octect[53]  = 00110101; //Value before code_group
    tx_octect[54]  = 00110110; //Value before code_group
    tx_octect[55]  = 00110111; //Value before code_group
    tx_octect[56]  = 00111000; //Value before code_group
    tx_octect[57]  = 00111001; //Value before code_group
    tx_octect[58]  = 00111010; //Value before code_group
    tx_octect[59]  = 00111011; //Value before code_group
    tx_octect[60]  = 00111100; //Value before code_group
    tx_octect[61]  = 00111101; //Value before code_group
    tx_octect[62]  = 00111110; //Value before code_group
    tx_octect[63]  = 00111111; //Value before code_group
    tx_octect[64]  = 01000000; //Value before code_group
    tx_octect[65]  = 01000001; //Value before code_group
    tx_octect[66]  = 01000010; //Value before code_group
    tx_octect[67]  = 01000011; //Value before code_group
    tx_octect[68]  = 01000100; //Value before code_group
    tx_octect[69]  = 01000101; //Value before code_group
    tx_octect[70]  = 01000110; //Value before code_group
    tx_octect[71]  = 01000111; //Value before code_group
    tx_octect[72]  = 01001000; //Value before code_group
    tx_octect[73]  = 01001001; //Value before code_group
    tx_octect[74]  = 01001010; //Value before code_group
    tx_octect[75]  = 01001011; //Value before code_group
    tx_octect[76]  = 01001100; //Value before code_group
    tx_octect[77]  = 01001101; //Value before code_group
    tx_octect[78]  = 01001110; //Value before code_group
    tx_octect[79]  = 01001111; //Value before code_group
    tx_octect[80]  = 01010000; //Value before code_group
    tx_octect[81]  = 01010001; //Value before code_group
    tx_octect[82]  = 01010010; //Value before code_group
    tx_octect[83]  = 01010011; //Value before code_group
    tx_octect[84]  = 01010100; //Value before code_group
    tx_octect[85]  = 01010101; //Value before code_group
    tx_octect[86]  = 01010110; //Value before code_group
    tx_octect[87]  = 01010111; //Value before code_group
    tx_octect[88]  = 01011000; //Value before code_group
    tx_octect[89]  = 01011001; //Value before code_group
    tx_octect[90]  = 01011010; //Value before code_group
    tx_octect[91]  = 01011011; //Value before code_group
    tx_octect[92]  = 01011100; //Value before code_group
    tx_octect[93]  = 01011101; //Value before code_group
    tx_octect[94]  = 01011110; //Value before code_group
    tx_octect[95]  = 01011111; //Value before code_group
    tx_octect[96]  = 01100000; //Value before code_group
    tx_octect[97]  = 01100001; //Value before code_group
    tx_octect[98]  = 01100010; //Value before code_group
    tx_octect[99]  = 01100011; //Value before code_group
    tx_octect[100] = 01100100; //Value before code_group
    tx_octect[101] = 01100101; //Value before code_group
    tx_octect[102] = 01100110; //Value before code_group
    tx_octect[103] = 01100111; //Value before code_group
    tx_octect[104] = 01101000; //Value before code_group
    tx_octect[105] = 01101001; //Value before code_group
    tx_octect[106] = 01101010; //Value before code_group
    tx_octect[107] = 01101011; //Value before code_group
    tx_octect[108] = 01101100; //Value before code_group
    tx_octect[109] = 01101101; //Value before code_group
    tx_octect[110] = 01101110; //Value before code_group
    tx_octect[111] = 01101111; //Value before code_group
    tx_octect[112] = 01110000; //Value before code_group
    tx_octect[113] = 01110001; //Value before code_group
    tx_octect[114] = 01110010; //Value before code_group
    tx_octect[115] = 01110011; //Value before code_group
    tx_octect[116] = 01110100; //Value before code_group
    tx_octect[117] = 01110101; //Value before code_group
    tx_octect[118] = 01110110; //Value before code_group
    tx_octect[119] = 01110111; //Value before code_group
    tx_octect[120] = 01111000; //Value before code_group
    tx_octect[121] = 01111001; //Value before code_group
    tx_octect[122] = 01111010; //Value before code_group
    tx_octect[123] = 01111011; //Value before code_group
    tx_octect[124] = 01111100; //Value before code_group
    tx_octect[125] = 01111101; //Value before code_group
    tx_octect[126] = 01111110; //Value before code_group
    tx_octect[127] = 01111111; //Value before code_group
    tx_octect[128] = 10000000; //Value before code_group
    tx_octect[129] = 10000001; //Value before code_group
    tx_octect[130] = 10000010; //Value before code_group
    tx_octect[131] = 10000011; //Value before code_group
    tx_octect[132] = 10000100; //Value before code_group
    tx_octect[133] = 10000101; //Value before code_group
    tx_octect[134] = 10000110; //Value before code_group
    tx_octect[135] = 10000111; //Value before code_group
    tx_octect[136] = 10001000; //Value before code_group
    tx_octect[137] = 10001001; //Value before code_group
    tx_octect[138] = 10001010; //Value before code_group
    tx_octect[139] = 10001011; //Value before code_group
    tx_octect[140] = 10001100; //Value before code_group
    tx_octect[141] = 10001101; //Value before code_group
    tx_octect[142] = 10001110; //Value before code_group
    tx_octect[143] = 10001111; //Value before code_group
    tx_octect[144] = 10010000; //Value before code_group
    tx_octect[145] = 10010001; //Value before code_group
    tx_octect[146] = 10010010; //Value before code_group
    tx_octect[147] = 10010011; //Value before code_group
    tx_octect[148] = 10010100; //Value before code_group
    tx_octect[149] = 10010101; //Value before code_group
    tx_octect[150] = 10010110; //Value before code_group
    tx_octect[151] = 10010111; //Value before code_group
    tx_octect[152] = 10011000; //Value before code_group
    tx_octect[153] = 10011001; //Value before code_group
    tx_octect[154] = 10011010; //Value before code_group
    tx_octect[155] = 10011011; //Value before code_group
    tx_octect[156] = 10011100; //Value before code_group
    tx_octect[157] = 10011101; //Value before code_group
    tx_octect[158] = 10011110; //Value before code_group
    tx_octect[159] = 10011111; //Value before code_group
    tx_octect[160] = 10100000; //Value before code_group
    tx_octect[161] = 10100001; //Value before code_group
    tx_octect[162] = 10100010; //Value before code_group
    tx_octect[163] = 10100011; //Value before code_group
    tx_octect[164] = 10100100; //Value before code_group
    tx_octect[165] = 10100101; //Value before code_group
    tx_octect[166] = 10100110; //Value before code_group
    tx_octect[167] = 10100111; //Value before code_group
    tx_octect[168] = 10101000; //Value before code_group
    tx_octect[169] = 10101001; //Value before code_group
    tx_octect[170] = 10101010; //Value before code_group
    tx_octect[171] = 10101011; //Value before code_group
    tx_octect[172] = 10101100; //Value before code_group
    tx_octect[173] = 10101101; //Value before code_group
    tx_octect[174] = 10101110; //Value before code_group
    tx_octect[175] = 10101111; //Value before code_group
    tx_octect[176] = 10110000; //Value before code_group
    tx_octect[177] = 10110001; //Value before code_group
    tx_octect[178] = 10110010; //Value before code_group
    tx_octect[179] = 10110011; //Value before code_group
    tx_octect[180] = 10110100; //Value before code_group
    tx_octect[181] = 10110101; //Value before code_group
    tx_octect[182] = 10110110; //Value before code_group
    tx_octect[183] = 10110111; //Value before code_group
    tx_octect[184] = 10111000; //Value before code_group
    tx_octect[185] = 10111001; //Value before code_group
    tx_octect[186] = 10111010; //Value before code_group
    tx_octect[187] = 10111011; //Value before code_group
    tx_octect[188] = 10111100; //Value before code_group
    tx_octect[189] = 10111101; //Value before code_group
    tx_octect[190] = 10111110; //Value before code_group
    tx_octect[191] = 10111111; //Value before code_group
    tx_octect[192] = 11000000; //Value before code_group
    tx_octect[193] = 11000001; //Value before code_group
    tx_octect[194] = 11000010; //Value before code_group
    tx_octect[195] = 11000011; //Value before code_group
    tx_octect[196] = 11000100; //Value before code_group
    tx_octect[197] = 11000101; //Value before code_group
    tx_octect[198] = 11000110; //Value before code_group
    tx_octect[199] = 11000111; //Value before code_group
    tx_octect[200] = 11001000; //Value before code_group
    tx_octect[201] = 11001001; //Value before code_group
    tx_octect[202] = 11001010; //Value before code_group
    tx_octect[203] = 11001011; //Value before code_group
    tx_octect[204] = 11001100; //Value before code_group
    tx_octect[205] = 11001101; //Value before code_group
    tx_octect[206] = 11001110; //Value before code_group
    tx_octect[207] = 11001111; //Value before code_group
    tx_octect[208] = 11010000; //Value before code_group
    tx_octect[209] = 11010001; //Value before code_group
    tx_octect[210] = 11010010; //Value before code_group
    tx_octect[211] = 11010011; //Value before code_group
    tx_octect[212] = 11010100; //Value before code_group
    tx_octect[213] = 11010101; //Value before code_group
    tx_octect[214] = 11010110; //Value before code_group
    tx_octect[215] = 11010111; //Value before code_group
    tx_octect[216] = 11011000; //Value before code_group
    tx_octect[217] = 11011001; //Value before code_group
    tx_octect[218] = 11011010; //Value before code_group
    tx_octect[219] = 11011011; //Value before code_group
    tx_octect[220] = 11011100; //Value before code_group
    tx_octect[221] = 11011101; //Value before code_group
    tx_octect[222] = 11011110; //Value before code_group
    tx_octect[223] = 11011111; //Value before code_group
    tx_octect[224] = 11100000; //Value before code_group
    tx_octect[225] = 11100001; //Value before code_group
    tx_octect[226] = 11100010; //Value before code_group
    tx_octect[227] = 11100011; //Value before code_group
    tx_octect[228] = 11100100; //Value before code_group
    tx_octect[229] = 11100101; //Value before code_group
    tx_octect[230] = 11100110; //Value before code_group
    tx_octect[231] = 11100111; //Value before code_group
    tx_octect[232] = 11101000; //Value before code_group
    tx_octect[233] = 11101001; //Value before code_group
    tx_octect[234] = 11101010; //Value before code_group
    tx_octect[235] = 11101011; //Value before code_group
    tx_octect[236] = 11101100; //Value before code_group
    tx_octect[237] = 11101101; //Value before code_group
    tx_octect[238] = 11101110; //Value before code_group
    tx_octect[239] = 11101111; //Value before code_group
    tx_octect[240] = 11110000; //Value before code_group
    tx_octect[241] = 11110001; //Value before code_group
    tx_octect[242] = 11110010; //Value before code_group
    tx_octect[243] = 11110011; //Value before code_group
    tx_octect[244] = 11110100; //Value before code_group
    tx_octect[245] = 11110101; //Value before code_group
    tx_octect[246] = 11110110; //Value before code_group
    tx_octect[247] = 11110111; //Value before code_group
    tx_octect[248] = 11111000; //Value before code_group
    tx_octect[249] = 11111001; //Value before code_group
    tx_octect[250] = 11111010; //Value before code_group
    tx_octect[251] = 11111011; //Value before code_group
    tx_octect[252] = 11111100; //Value before code_group
    tx_octect[253] = 11111101; //Value before code_group
    tx_octect[254] = 11111110; //Value before code_group
    tx_octect[255] = 11111111; //Value before code_group
    tx_octect[256] = 00011100; //Value before code_group
    tx_octect[257] = 00111100; //Value before code_group
    tx_octect[258] = 01011100; //Value before code_group
    tx_octect[259] = 01111100; //Value before code_group
    tx_octect[260] = 10011100; //Value before code_group
    tx_octect[261] = 10111100; //Value before code_group
    tx_octect[262] = 11011100; //Value before code_group
    tx_octect[263] = 11111100; //Value before code_group
    tx_octect[264] = 11110111; //Value before code_group
    tx_octect[265] = 11111011; //Value before code_group
    tx_octect[266] = 11111101; //Value before code_group
    tx_octect[267] = 11111110; //Value before code_group
    
    
                                           //Impares
    code_group_Imp[0]   = 10'b1001110100; //Octect Value in Binary: 000 00000
    code_group_Imp[1]   = 10'b0111010100; //Octect Value in Binary: 000 00001
    code_group_Imp[2]   = 10'b1011010100; //Octect Value in Binary: 000 00010
    code_group_Imp[3]   = 10'b1100011011; //Octect Value in Binary: 000 00011
    code_group_Imp[4]   = 10'b1101010100; //Octect Value in Binary: 000 00100
    code_group_Imp[5]   = 10'b1010011011; //Octect Value in Binary: 000 00101
    code_group_Imp[6]   = 10'b0110011011; //Octect Value in Binary: 000 00110
    code_group_Imp[7]   = 10'b1110001011; //Octect Value in Binary: 000 00111
    code_group_Imp[8]   = 10'b1110010100; //Octect Value in Binary: 000 01000
    code_group_Imp[9]   = 10'b1001011011; //Octect Value in Binary: 000 01001
    code_group_Imp[10]  = 10'b0101011011; //Octect Value in Binary: 000 01010
    code_group_Imp[11]  = 10'b1101001011; //Octect Value in Binary: 000 01011
    code_group_Imp[12]  = 10'b0011011011; //Octect Value in Binary: 000 01100
    code_group_Imp[13]  = 10'b1011001011; //Octect Value in Binary: 000 01101
    code_group_Imp[14]  = 10'b0111001011; //Octect Value in Binary: 000 01110
    code_group_Imp[15]  = 10'b0101110100; //Octect Value in Binary: 000 01111
    code_group_Imp[16]  = 10'b0110110100; //Octect Value in Binary: 000 10000
    code_group_Imp[17]  = 10'b1000111011; //Octect Value in Binary: 000 10001
    code_group_Imp[18]  = 10'b0100111011; //Octect Value in Binary: 000 10010
    code_group_Imp[19]  = 10'b1100101011; //Octect Value in Binary: 000 10011
    code_group_Imp[20]  = 10'b0010111011; //Octect Value in Binary: 000 10100
    code_group_Imp[21]  = 10'b1010101011; //Octect Value in Binary: 000 10101
    code_group_Imp[22]  = 10'b0110101011; //Octect Value in Binary: 000 10110
    code_group_Imp[23]  = 10'b1110100100; //Octect Value in Binary: 000 10111
    code_group_Imp[24]  = 10'b1100110100; //Octect Value in Binary: 000 11000
    code_group_Imp[25]  = 10'b1001101011; //Octect Value in Binary: 000 11001
    code_group_Imp[26]  = 10'b0101101011; //Octect Value in Binary: 000 11010
    code_group_Imp[27]  = 10'b1101100100; //Octect Value in Binary: 000 11011
    code_group_Imp[28]  = 10'b0011101011; //Octect Value in Binary: 000 11100
    code_group_Imp[29]  = 10'b1011100100; //Octect Value in Binary: 000 11101
    code_group_Imp[30]  = 10'b0111100100; //Octect Value in Binary: 000 11110
    code_group_Imp[31]  = 10'b1010110100; //Octect Value in Binary: 000 11111
    code_group_Imp[32]  = 10'b1001111001; //Octect Value in Binary: 001 00000
    code_group_Imp[33]  = 10'b0111011001; //Octect Value in Binary: 001 00001
    code_group_Imp[34]  = 10'b1011011001; //Octect Value in Binary: 001 00010
    code_group_Imp[35]  = 10'b1100011001; //Octect Value in Binary: 001 00011
    code_group_Imp[36]  = 10'b1101011001; //Octect Value in Binary: 001 00100
    code_group_Imp[37]  = 10'b1010011001; //Octect Value in Binary: 001 00101
    code_group_Imp[38]  = 10'b0110011001; //Octect Value in Binary: 001 00110
    code_group_Imp[39]  = 10'b1110001001; //Octect Value in Binary: 001 00111
    code_group_Imp[40]  = 10'b1110011001; //Octect Value in Binary: 001 01000
    code_group_Imp[41]  = 10'b1001011001; //Octect Value in Binary: 001 01001
    code_group_Imp[42]  = 10'b0101011001; //Octect Value in Binary: 001 01010
    code_group_Imp[43]  = 10'b1101001001; //Octect Value in Binary: 001 01011
    code_group_Imp[44]  = 10'b0011011001; //Octect Value in Binary: 001 01100
    code_group_Imp[45]  = 10'b1011001001; //Octect Value in Binary: 001 01101
    code_group_Imp[46]  = 10'b0111001001; //Octect Value in Binary: 001 01110
    code_group_Imp[47]  = 10'b0101111001; //Octect Value in Binary: 001 01111
    code_group_Imp[48]  = 10'b0110111001; //Octect Value in Binary: 001 10000
    code_group_Imp[49]  = 10'b1000111001; //Octect Value in Binary: 001 10001
    code_group_Imp[50]  = 10'b0100111001; //Octect Value in Binary: 001 10010
    code_group_Imp[51]  = 10'b1100101001; //Octect Value in Binary: 001 10011
    code_group_Imp[52]  = 10'b0010111001; //Octect Value in Binary: 001 10100
    code_group_Imp[53]  = 10'b1010101001; //Octect Value in Binary: 001 10101
    code_group_Imp[54]  = 10'b0110101001; //Octect Value in Binary: 001 10110
    code_group_Imp[55]  = 10'b1110101001; //Octect Value in Binary: 001 10111
    code_group_Imp[56]  = 10'b1100111001; //Octect Value in Binary: 001 11000
    code_group_Imp[57]  = 10'b1001101001; //Octect Value in Binary: 001 11001
    code_group_Imp[58]  = 10'b0101101001; //Octect Value in Binary: 001 11010
    code_group_Imp[59]  = 10'b1101101001; //Octect Value in Binary: 001 11011
    code_group_Imp[60]  = 10'b0011101001; //Octect Value in Binary: 001 11100
    code_group_Imp[61]  = 10'b1011101001; //Octect Value in Binary: 001 11101
    code_group_Imp[62]  = 10'b0111101001; //Octect Value in Binary: 001 11110
    code_group_Imp[63]  = 10'b1010111001; //Octect Value in Binary: 001 11111
    code_group_Imp[64]  = 10'b1001110101; //Octect Value in Binary: 010 00000
    code_group_Imp[65]  = 10'b0111010101; //Octect Value in Binary: 010 00001
    code_group_Imp[66]  = 10'b1011010101; //Octect Value in Binary: 010 00010
    code_group_Imp[67]  = 10'b1100010101; //Octect Value in Binary: 010 00011
    code_group_Imp[68]  = 10'b1101010101; //Octect Value in Binary: 010 00100
    code_group_Imp[69]  = 10'b1010010101; //Octect Value in Binary: 010 00101
    code_group_Imp[70]  = 10'b0110010101; //Octect Value in Binary: 010 00110
    code_group_Imp[71]  = 10'b1110000101; //Octect Value in Binary: 010 00111
    code_group_Imp[72]  = 10'b1110010101; //Octect Value in Binary: 010 01000
    code_group_Imp[73]  = 10'b1001010101; //Octect Value in Binary: 010 01001
    code_group_Imp[74]  = 10'b0101010101; //Octect Value in Binary: 010 01010
    code_group_Imp[75]  = 10'b1101000101; //Octect Value in Binary: 010 01011
    code_group_Imp[76]  = 10'b0011010101; //Octect Value in Binary: 010 01100
    code_group_Imp[77]  = 10'b1011000101; //Octect Value in Binary: 010 01101
    code_group_Imp[78]  = 10'b0111000101; //Octect Value in Binary: 010 01110
    code_group_Imp[79]  = 10'b0101110101; //Octect Value in Binary: 010 01111
    code_group_Imp[80]  = 10'b0110110101; //Octect Value in Binary: 010 10000
    code_group_Imp[81]  = 10'b1000110101; //Octect Value in Binary: 010 10001
    code_group_Imp[82]  = 10'b0100110101; //Octect Value in Binary: 010 10010
    code_group_Imp[83]  = 10'b1100100101; //Octect Value in Binary: 010 10011
    code_group_Imp[84]  = 10'b0010110101; //Octect Value in Binary: 010 10100
    code_group_Imp[85]  = 10'b1010100101; //Octect Value in Binary: 010 10101
    code_group_Imp[86]  = 10'b0110100101; //Octect Value in Binary: 010 10110
    code_group_Imp[87]  = 10'b1110100101; //Octect Value in Binary: 010 10111
    code_group_Imp[88]  = 10'b1100110101; //Octect Value in Binary: 010 11000
    code_group_Imp[89]  = 10'b1001100101; //Octect Value in Binary: 010 11001
    code_group_Imp[90]  = 10'b0101100101; //Octect Value in Binary: 010 11010
    code_group_Imp[91]  = 10'b1101100101; //Octect Value in Binary: 010 11011
    code_group_Imp[92]  = 10'b0011100101; //Octect Value in Binary: 010 11100
    code_group_Imp[93]  = 10'b1011100101; //Octect Value in Binary: 010 11101
    code_group_Imp[94]  = 10'b0111100101; //Octect Value in Binary: 010 11110
    code_group_Imp[95]  = 10'b1010110101; //Octect Value in Binary: 010 11111
    code_group_Imp[96]  = 10'b1001110011; //Octect Value in Binary: 011 00000
    code_group_Imp[97]  = 10'b0111010011; //Octect Value in Binary: 011 00001
    code_group_Imp[98]  = 10'b1011010011; //Octect Value in Binary: 011 00010
    code_group_Imp[99]  = 10'b1100011100; //Octect Value in Binary: 011 00011
    code_group_Imp[100] = 10'b1101010011; //Octect Value in Binary: 011 00100
    code_group_Imp[101] = 10'b1010011100; //Octect Value in Binary: 011 00101
    code_group_Imp[102] = 10'b0110011100; //Octect Value in Binary: 011 00110
    code_group_Imp[103] = 10'b1110001100; //Octect Value in Binary: 011 00111
    code_group_Imp[104] = 10'b1110010011; //Octect Value in Binary: 011 01000
    code_group_Imp[105] = 10'b1001011100; //Octect Value in Binary: 011 01001
    code_group_Imp[106] = 10'b0101011100; //Octect Value in Binary: 011 01010
    code_group_Imp[107] = 10'b1101001100; //Octect Value in Binary: 011 01011
    code_group_Imp[108] = 10'b0011011100; //Octect Value in Binary: 011 01100
    code_group_Imp[109] = 10'b1011001100; //Octect Value in Binary: 011 01101
    code_group_Imp[110] = 10'b0111001100; //Octect Value in Binary: 011 01110
    code_group_Imp[111] = 10'b0101110011; //Octect Value in Binary: 011 01111
    code_group_Imp[112] = 10'b0110110011; //Octect Value in Binary: 011 10000
    code_group_Imp[113] = 10'b1000111100; //Octect Value in Binary: 011 10001
    code_group_Imp[114] = 10'b0100111100; //Octect Value in Binary: 011 10010
    code_group_Imp[115] = 10'b1100101100; //Octect Value in Binary: 011 10011
    code_group_Imp[116] = 10'b0010111100; //Octect Value in Binary: 011 10100
    code_group_Imp[117] = 10'b1010101100; //Octect Value in Binary: 011 10101
    code_group_Imp[118] = 10'b0110101100; //Octect Value in Binary: 011 10110
    code_group_Imp[119] = 10'b1110100011; //Octect Value in Binary: 011 10111
    code_group_Imp[120] = 10'b1100110011; //Octect Value in Binary: 011 11000
    code_group_Imp[121] = 10'b1001101100; //Octect Value in Binary: 011 11001
    code_group_Imp[122] = 10'b0101101100; //Octect Value in Binary: 011 11010
    code_group_Imp[123] = 10'b1101100011; //Octect Value in Binary: 011 11011
    code_group_Imp[124] = 10'b0011101100; //Octect Value in Binary: 011 11100
    code_group_Imp[125] = 10'b1011100011; //Octect Value in Binary: 011 11101
    code_group_Imp[126] = 10'b0111100011; //Octect Value in Binary: 011 11110
    code_group_Imp[127] = 10'b1010110011; //Octect Value in Binary: 011 11111
    code_group_Imp[128] = 10'b1001110010; //Octect Value in Binary: 100 00000
    code_group_Imp[129] = 10'b0111010010; //Octect Value in Binary: 100 00001
    code_group_Imp[130] = 10'b1011010010; //Octect Value in Binary: 100 00010
    code_group_Imp[131] = 10'b1100011101; //Octect Value in Binary: 100 00011
    code_group_Imp[132] = 10'b1101010010; //Octect Value in Binary: 100 00100
    code_group_Imp[133] = 10'b1010011101; //Octect Value in Binary: 100 00101
    code_group_Imp[134] = 10'b0110011101; //Octect Value in Binary: 100 00110
    code_group_Imp[135] = 10'b1110001101; //Octect Value in Binary: 100 00111
    code_group_Imp[136] = 10'b1110010010; //Octect Value in Binary: 100 01000
    code_group_Imp[137] = 10'b1001011101; //Octect Value in Binary: 100 01001
    code_group_Imp[138] = 10'b0101011101; //Octect Value in Binary: 100 01010
    code_group_Imp[139] = 10'b1101001101; //Octect Value in Binary: 100 01011
    code_group_Imp[140] = 10'b0011011101; //Octect Value in Binary: 100 01100
    code_group_Imp[141] = 10'b1011001101; //Octect Value in Binary: 100 01101
    code_group_Imp[142] = 10'b0111001101; //Octect Value in Binary: 100 01110
    code_group_Imp[143] = 10'b0101110010; //Octect Value in Binary: 100 01111
    code_group_Imp[144] = 10'b0110110010; //Octect Value in Binary: 100 10000
    code_group_Imp[145] = 10'b1000111101; //Octect Value in Binary: 100 10001
    code_group_Imp[146] = 10'b0100111101; //Octect Value in Binary: 100 10010
    code_group_Imp[147] = 10'b1100101101; //Octect Value in Binary: 100 10011
    code_group_Imp[148] = 10'b0010111101; //Octect Value in Binary: 100 10100
    code_group_Imp[149] = 10'b1010101101; //Octect Value in Binary: 100 10101
    code_group_Imp[150] = 10'b0110101101; //Octect Value in Binary: 100 10110
    code_group_Imp[151] = 10'b1110100010; //Octect Value in Binary: 100 10111
    code_group_Imp[152] = 10'b1100110010; //Octect Value in Binary: 100 11000
    code_group_Imp[153] = 10'b1001101101; //Octect Value in Binary: 100 11001
    code_group_Imp[154] = 10'b0101101101; //Octect Value in Binary: 100 11010
    code_group_Imp[155] = 10'b1101100010; //Octect Value in Binary: 100 11011
    code_group_Imp[156] = 10'b0011101101; //Octect Value in Binary: 100 11100
    code_group_Imp[157] = 10'b1011100010; //Octect Value in Binary: 100 11101
    code_group_Imp[158] = 10'b0111100010; //Octect Value in Binary: 100 11110
    code_group_Imp[159] = 10'b1010110010; //Octect Value in Binary: 100 11111
    code_group_Imp[160] = 10'b1001111010; //Octect Value in Binary: 101 00000
    code_group_Imp[161] = 10'b0111011010; //Octect Value in Binary: 101 00001
    code_group_Imp[162] = 10'b1011011010; //Octect Value in Binary: 101 00010
    code_group_Imp[163] = 10'b1100011010; //Octect Value in Binary: 101 00011
    code_group_Imp[164] = 10'b1101011010; //Octect Value in Binary: 101 00100
    code_group_Imp[165] = 10'b1010011010; //Octect Value in Binary: 101 00101
    code_group_Imp[166] = 10'b0110011010; //Octect Value in Binary: 101 00110
    code_group_Imp[167] = 10'b1110001010; //Octect Value in Binary: 101 00111
    code_group_Imp[168] = 10'b1110011010; //Octect Value in Binary: 101 01000
    code_group_Imp[169] = 10'b1001011010; //Octect Value in Binary: 101 01001
    code_group_Imp[170] = 10'b0101011010; //Octect Value in Binary: 101 01010
    code_group_Imp[171] = 10'b1101001010; //Octect Value in Binary: 101 01011
    code_group_Imp[172] = 10'b0011011010; //Octect Value in Binary: 101 01100
    code_group_Imp[173] = 10'b1011001010; //Octect Value in Binary: 101 01101
    code_group_Imp[174] = 10'b0111001010; //Octect Value in Binary: 101 01110
    code_group_Imp[175] = 10'b0101111010; //Octect Value in Binary: 101 01111
    code_group_Imp[176] = 10'b0110111010; //Octect Value in Binary: 101 10000
    code_group_Imp[177] = 10'b1000111010; //Octect Value in Binary: 101 10001
    code_group_Imp[178] = 10'b0100111010; //Octect Value in Binary: 101 10010
    code_group_Imp[179] = 10'b1100101010; //Octect Value in Binary: 101 10011
    code_group_Imp[180] = 10'b0010111010; //Octect Value in Binary: 101 10100
    code_group_Imp[181] = 10'b1010101010; //Octect Value in Binary: 101 10101
    code_group_Imp[182] = 10'b0110101010; //Octect Value in Binary: 101 10110
    code_group_Imp[183] = 10'b1110101010; //Octect Value in Binary: 101 10111
    code_group_Imp[184] = 10'b1100111010; //Octect Value in Binary: 101 11000
    code_group_Imp[185] = 10'b1001101010; //Octect Value in Binary: 101 11001
    code_group_Imp[186] = 10'b0101101010; //Octect Value in Binary: 101 11010
    code_group_Imp[187] = 10'b1101101010; //Octect Value in Binary: 101 11011
    code_group_Imp[188] = 10'b0011101010; //Octect Value in Binary: 101 11100
    code_group_Imp[189] = 10'b1011101010; //Octect Value in Binary: 101 11101
    code_group_Imp[190] = 10'b0111101010; //Octect Value in Binary: 101 11110
    code_group_Imp[191] = 10'b1010111010; //Octect Value in Binary: 101 11111
    code_group_Imp[192] = 10'b1001110110; //Octect Value in Binary: 110 00000
    code_group_Imp[193] = 10'b0111010110; //Octect Value in Binary: 110 00001
    code_group_Imp[194] = 10'b1011010110; //Octect Value in Binary: 110 00010
    code_group_Imp[195] = 10'b1100010110; //Octect Value in Binary: 110 00011
    code_group_Imp[196] = 10'b1101010110; //Octect Value in Binary: 110 00100
    code_group_Imp[197] = 10'b1010010110; //Octect Value in Binary: 110 00101
    code_group_Imp[198] = 10'b0110010110; //Octect Value in Binary: 110 00110
    code_group_Imp[199] = 10'b1110000110; //Octect Value in Binary: 110 00111
    code_group_Imp[200] = 10'b1110010110; //Octect Value in Binary: 110 01000
    code_group_Imp[201] = 10'b1001010110; //Octect Value in Binary: 110 01001
    code_group_Imp[202] = 10'b0101010110; //Octect Value in Binary: 110 01010
    code_group_Imp[203] = 10'b1101000110; //Octect Value in Binary: 110 01011
    code_group_Imp[204] = 10'b0011010110; //Octect Value in Binary: 110 01100
    code_group_Imp[205] = 10'b1011000110; //Octect Value in Binary: 110 01101
    code_group_Imp[206] = 10'b0111000110; //Octect Value in Binary: 110 01110
    code_group_Imp[207] = 10'b0101110110; //Octect Value in Binary: 110 01111
    code_group_Imp[208] = 10'b0110110110; //Octect Value in Binary: 110 10000
    code_group_Imp[209] = 10'b1000110110; //Octect Value in Binary: 110 10001
    code_group_Imp[210] = 10'b0100110110; //Octect Value in Binary: 110 10010
    code_group_Imp[211] = 10'b1100100110; //Octect Value in Binary: 110 10011
    code_group_Imp[212] = 10'b0010110110; //Octect Value in Binary: 110 10100
    code_group_Imp[213] = 10'b1010100110; //Octect Value in Binary: 110 10101
    code_group_Imp[214] = 10'b0110100110; //Octect Value in Binary: 110 10110
    code_group_Imp[215] = 10'b1110100110; //Octect Value in Binary: 110 10111
    code_group_Imp[216] = 10'b1100110110; //Octect Value in Binary: 110 11000
    code_group_Imp[217] = 10'b1001100110; //Octect Value in Binary: 110 11001
    code_group_Imp[218] = 10'b0101100110; //Octect Value in Binary: 110 11010
    code_group_Imp[219] = 10'b1101100110; //Octect Value in Binary: 110 11011
    code_group_Imp[220] = 10'b0011100110; //Octect Value in Binary: 110 11100
    code_group_Imp[221] = 10'b1011100110; //Octect Value in Binary: 110 11101
    code_group_Imp[222] = 10'b0111100110; //Octect Value in Binary: 110 11110
    code_group_Imp[223] = 10'b1010110110; //Octect Value in Binary: 110 11111
    code_group_Imp[224] = 10'b1001110001; //Octect Value in Binary: 111 00000
    code_group_Imp[225] = 10'b0111010001; //Octect Value in Binary: 111 00001
    code_group_Imp[226] = 10'b1011010001; //Octect Value in Binary: 111 00010
    code_group_Imp[227] = 10'b1100011110; //Octect Value in Binary: 111 00011
    code_group_Imp[228] = 10'b1101010001; //Octect Value in Binary: 111 00100
    code_group_Imp[229] = 10'b1010011110; //Octect Value in Binary: 111 00101
    code_group_Imp[230] = 10'b0110011110; //Octect Value in Binary: 111 00110
    code_group_Imp[231] = 10'b1110001110; //Octect Value in Binary: 111 00111
    code_group_Imp[232] = 10'b1110010001; //Octect Value in Binary: 111 01000
    code_group_Imp[233] = 10'b1001011110; //Octect Value in Binary: 111 01001
    code_group_Imp[234] = 10'b0101011110; //Octect Value in Binary: 111 01010
    code_group_Imp[235] = 10'b1101001110; //Octect Value in Binary: 111 01011
    code_group_Imp[236] = 10'b0011011110; //Octect Value in Binary: 111 01100
    code_group_Imp[237] = 10'b1011001110; //Octect Value in Binary: 111 01101
    code_group_Imp[238] = 10'b0111001110; //Octect Value in Binary: 111 01110
    code_group_Imp[239] = 10'b0101110001; //Octect Value in Binary: 111 01111
    code_group_Imp[240] = 10'b0110110001; //Octect Value in Binary: 111 10000
    code_group_Imp[241] = 10'b1000110111; //Octect Value in Binary: 111 10001
    code_group_Imp[242] = 10'b0100110111; //Octect Value in Binary: 111 10010
    code_group_Imp[243] = 10'b1100101110; //Octect Value in Binary: 111 10011
    code_group_Imp[244] = 10'b0010110111; //Octect Value in Binary: 111 10100
    code_group_Imp[245] = 10'b1010101110; //Octect Value in Binary: 111 10101
    code_group_Imp[246] = 10'b0110101110; //Octect Value in Binary: 111 10110
    code_group_Imp[247] = 10'b1110100001; //Octect Value in Binary: 111 10111
    code_group_Imp[248] = 10'b1100110001; //Octect Value in Binary: 111 11000
    code_group_Imp[249] = 10'b1001101110; //Octect Value in Binary: 111 11001
    code_group_Imp[250] = 10'b0101101110; //Octect Value in Binary: 111 11010
    code_group_Imp[251] = 10'b1101100001; //Octect Value in Binary: 111 11011
    code_group_Imp[252] = 10'b0011101110; //Octect Value in Binary: 111 11100
    code_group_Imp[253] = 10'b1011100001; //Octect Value in Binary: 111 11101
    code_group_Imp[254] = 10'b0111100001; //Octect Value in Binary: 111 11110
    code_group_Imp[255] = 10'b1010110001; //Octect Value in Binary: 111 11111
    code_group_Imp[256] = 10'b0011110100; //Octect Value in Binary: 000 11100
    code_group_Imp[257] = 10'b0011111001; //Octect Value in Binary: 001 11100
    code_group_Imp[258] = 10'b0011110101; //Octect Value in Binary: 010 11100
    code_group_Imp[259] = 10'b0011110011; //Octect Value in Binary: 011 11100
    code_group_Imp[260] = 10'b0011110010; //Octect Value in Binary: 100 11100
    code_group_Imp[261] = 10'b0011111010; //Octect Value in Binary: 101 11100
    code_group_Imp[262] = 10'b0011110110; //Octect Value in Binary: 110 11100
    code_group_Imp[263] = 10'b0011111000; //Octect Value in Binary: 111 11100
    code_group_Imp[264] = 10'b1110101000; //Octect Value in Binary: 111 10111
    code_group_Imp[265] = 10'b1101101000; //Octect Value in Binary: 111 11011
    code_group_Imp[266] = 10'b1011101000; //Octect Value in Binary: 111 11101
    code_group_Imp[267] = 10'b0111101000; //Octect Value in Binary: 111 11110
    
                                           //Pares
    code_group_Par[0]   = 10'b0110001011; //Octect Value in Binary: 000 00000
    code_group_Par[1]   = 10'b1000101011; //Octect Value in Binary: 000 00001
    code_group_Par[2]   = 10'b0100101011; //Octect Value in Binary: 000 00010
    code_group_Par[3]   = 10'b1100010100; //Octect Value in Binary: 000 00011
    code_group_Par[4]   = 10'b0010101011; //Octect Value in Binary: 000 00100
    code_group_Par[5]   = 10'b1010010100; //Octect Value in Binary: 000 00101
    code_group_Par[6]   = 10'b0110010100; //Octect Value in Binary: 000 00110
    code_group_Par[7]   = 10'b0001110100; //Octect Value in Binary: 000 00111
    code_group_Par[8]   = 10'b0001101011; //Octect Value in Binary: 000 01000
    code_group_Par[9]   = 10'b1001010100; //Octect Value in Binary: 000 01001
    code_group_Par[10]  = 10'b0101010100; //Octect Value in Binary: 000 01010
    code_group_Par[11]  = 10'b1101000100; //Octect Value in Binary: 000 01011
    code_group_Par[12]  = 10'b0011010100; //Octect Value in Binary: 000 01100
    code_group_Par[13]  = 10'b1011000100; //Octect Value in Binary: 000 01101
    code_group_Par[14]  = 10'b0111000100; //Octect Value in Binary: 000 01110
    code_group_Par[15]  = 10'b1010001011; //Octect Value in Binary: 000 01111
    code_group_Par[16]  = 10'b1001001011; //Octect Value in Binary: 000 10000
    code_group_Par[17]  = 10'b1000110100; //Octect Value in Binary: 000 10001
    code_group_Par[18]  = 10'b0100110100; //Octect Value in Binary: 000 10010
    code_group_Par[19]  = 10'b1100100100; //Octect Value in Binary: 000 10011
    code_group_Par[20]  = 10'b0010110100; //Octect Value in Binary: 000 10100
    code_group_Par[21]  = 10'b1010100100; //Octect Value in Binary: 000 10101
    code_group_Par[22]  = 10'b0110100100; //Octect Value in Binary: 000 10110
    code_group_Par[23]  = 10'b0001011011; //Octect Value in Binary: 000 10111
    code_group_Par[24]  = 10'b0011001011; //Octect Value in Binary: 000 11000
    code_group_Par[25]  = 10'b1001100100; //Octect Value in Binary: 000 11001
    code_group_Par[26]  = 10'b0101100100; //Octect Value in Binary: 000 11010
    code_group_Par[27]  = 10'b0010011011; //Octect Value in Binary: 000 11011
    code_group_Par[28]  = 10'b0011100100; //Octect Value in Binary: 000 11100
    code_group_Par[29]  = 10'b0100011011; //Octect Value in Binary: 000 11101
    code_group_Par[30]  = 10'b1000011011; //Octect Value in Binary: 000 11110
    code_group_Par[31]  = 10'b0101001011; //Octect Value in Binary: 000 11111
    code_group_Par[32]  = 10'b0110001001; //Octect Value in Binary: 001 00000
    code_group_Par[33]  = 10'b1000101001; //Octect Value in Binary: 001 00001
    code_group_Par[34]  = 10'b0100101001; //Octect Value in Binary: 001 00010
    code_group_Par[35]  = 10'b1100011001; //Octect Value in Binary: 001 00011
    code_group_Par[36]  = 10'b0010101001; //Octect Value in Binary: 001 00100
    code_group_Par[37]  = 10'b1010011001; //Octect Value in Binary: 001 00101
    code_group_Par[38]  = 10'b0110011001; //Octect Value in Binary: 001 00110
    code_group_Par[39]  = 10'b0001111001; //Octect Value in Binary: 001 00111
    code_group_Par[40]  = 10'b0001101001; //Octect Value in Binary: 001 01000
    code_group_Par[41]  = 10'b1001011001; //Octect Value in Binary: 001 01001
    code_group_Par[42]  = 10'b0101011001; //Octect Value in Binary: 001 01010
    code_group_Par[43]  = 10'b1101001001; //Octect Value in Binary: 001 01011
    code_group_Par[44]  = 10'b0011011001; //Octect Value in Binary: 001 01100
    code_group_Par[45]  = 10'b1011001001; //Octect Value in Binary: 001 01101
    code_group_Par[46]  = 10'b0111001001; //Octect Value in Binary: 001 01110
    code_group_Par[47]  = 10'b1010001001; //Octect Value in Binary: 001 01111
    code_group_Par[48]  = 10'b1001001001; //Octect Value in Binary: 001 10000
    code_group_Par[49]  = 10'b1000111001; //Octect Value in Binary: 001 10001
    code_group_Par[50]  = 10'b0100111001; //Octect Value in Binary: 001 10010
    code_group_Par[51]  = 10'b1100101001; //Octect Value in Binary: 001 10011
    code_group_Par[52]  = 10'b0010111001; //Octect Value in Binary: 001 10100
    code_group_Par[53]  = 10'b1010101001; //Octect Value in Binary: 001 10101
    code_group_Par[54]  = 10'b0110101001; //Octect Value in Binary: 001 10110
    code_group_Par[55]  = 10'b0001011001; //Octect Value in Binary: 001 10111
    code_group_Par[56]  = 10'b0011001001; //Octect Value in Binary: 001 11000
    code_group_Par[57]  = 10'b1001101001; //Octect Value in Binary: 001 11001
    code_group_Par[58]  = 10'b0101101001; //Octect Value in Binary: 001 11010
    code_group_Par[59]  = 10'b0010011001; //Octect Value in Binary: 001 11011
    code_group_Par[60]  = 10'b0011101001; //Octect Value in Binary: 001 11100
    code_group_Par[61]  = 10'b0100011001; //Octect Value in Binary: 001 11101
    code_group_Par[62]  = 10'b1000011001; //Octect Value in Binary: 001 11110
    code_group_Par[63]  = 10'b0101001001; //Octect Value in Binary: 001 11111
    code_group_Par[64]  = 10'b0110000101; //Octect Value in Binary: 010 00000
    code_group_Par[65]  = 10'b1000100101; //Octect Value in Binary: 010 00001
    code_group_Par[66]  = 10'b0100100101; //Octect Value in Binary: 010 00010
    code_group_Par[67]  = 10'b1100010101; //Octect Value in Binary: 010 00011
    code_group_Par[68]  = 10'b0010100101; //Octect Value in Binary: 010 00100
    code_group_Par[69]  = 10'b1010010101; //Octect Value in Binary: 010 00101
    code_group_Par[70]  = 10'b0110010101; //Octect Value in Binary: 010 00110
    code_group_Par[71]  = 10'b0001110101; //Octect Value in Binary: 010 00111
    code_group_Par[72]  = 10'b0001100101; //Octect Value in Binary: 010 01000
    code_group_Par[73]  = 10'b1001010101; //Octect Value in Binary: 010 01001
    code_group_Par[74]  = 10'b0101010101; //Octect Value in Binary: 010 01010
    code_group_Par[75]  = 10'b1101000101; //Octect Value in Binary: 010 01011
    code_group_Par[76]  = 10'b0011010101; //Octect Value in Binary: 010 01100
    code_group_Par[77]  = 10'b1011000101; //Octect Value in Binary: 010 01101
    code_group_Par[78]  = 10'b0111000101; //Octect Value in Binary: 010 01110
    code_group_Par[79]  = 10'b1010000101; //Octect Value in Binary: 010 01111
    code_group_Par[80]  = 10'b1001000101; //Octect Value in Binary: 010 10000
    code_group_Par[81]  = 10'b1000110101; //Octect Value in Binary: 010 10001
    code_group_Par[82]  = 10'b0100110101; //Octect Value in Binary: 010 10010
    code_group_Par[83]  = 10'b1100100101; //Octect Value in Binary: 010 10011
    code_group_Par[84]  = 10'b0010110101; //Octect Value in Binary: 010 10100
    code_group_Par[85]  = 10'b1010100101; //Octect Value in Binary: 010 10101
    code_group_Par[86]  = 10'b0110100101; //Octect Value in Binary: 010 10110
    code_group_Par[87]  = 10'b0001010101; //Octect Value in Binary: 010 10111
    code_group_Par[88]  = 10'b0011000101; //Octect Value in Binary: 010 11000
    code_group_Par[89]  = 10'b1001100101; //Octect Value in Binary: 010 11001
    code_group_Par[90]  = 10'b0101100101; //Octect Value in Binary: 010 11010
    code_group_Par[91]  = 10'b0010010101; //Octect Value in Binary: 010 11011
    code_group_Par[92]  = 10'b0011100101; //Octect Value in Binary: 010 11100
    code_group_Par[93]  = 10'b0100010101; //Octect Value in Binary: 010 11101
    code_group_Par[94]  = 10'b1000010101; //Octect Value in Binary: 010 11110
    code_group_Par[95]  = 10'b0101000101; //Octect Value in Binary: 010 11111
    code_group_Par[96]  = 10'b0110001100; //Octect Value in Binary: 011 00000
    code_group_Par[97]  = 10'b1000101100; //Octect Value in Binary: 011 00001
    code_group_Par[98]  = 10'b0100101100; //Octect Value in Binary: 011 00010
    code_group_Par[99]  = 10'b1100010011; //Octect Value in Binary: 011 00011
    code_group_Par[100] = 10'b0010101100; //Octect Value in Binary: 011 00100
    code_group_Par[101] = 10'b1010010011; //Octect Value in Binary: 011 00101
    code_group_Par[102] = 10'b0110010011; //Octect Value in Binary: 011 00110
    code_group_Par[103] = 10'b0001110011; //Octect Value in Binary: 011 00111
    code_group_Par[104] = 10'b0001101100; //Octect Value in Binary: 011 01000
    code_group_Par[105] = 10'b1001010011; //Octect Value in Binary: 011 01001
    code_group_Par[106] = 10'b0101010011; //Octect Value in Binary: 011 01010
    code_group_Par[107] = 10'b1101000011; //Octect Value in Binary: 011 01011
    code_group_Par[108] = 10'b0011010011; //Octect Value in Binary: 011 01100
    code_group_Par[109] = 10'b1011000011; //Octect Value in Binary: 011 01101
    code_group_Par[110] = 10'b0111000011; //Octect Value in Binary: 011 01110
    code_group_Par[111] = 10'b1010001100; //Octect Value in Binary: 011 01111
    code_group_Par[112] = 10'b1001001100; //Octect Value in Binary: 011 10000
    code_group_Par[113] = 10'b1000110011; //Octect Value in Binary: 011 10001
    code_group_Par[114] = 10'b0100110011; //Octect Value in Binary: 011 10010
    code_group_Par[115] = 10'b1100100011; //Octect Value in Binary: 011 10011
    code_group_Par[116] = 10'b0010110011; //Octect Value in Binary: 011 10100
    code_group_Par[117] = 10'b1010100011; //Octect Value in Binary: 011 10101
    code_group_Par[118] = 10'b0110100011; //Octect Value in Binary: 011 10110
    code_group_Par[119] = 10'b0001011100; //Octect Value in Binary: 011 10111
    code_group_Par[120] = 10'b0011001100; //Octect Value in Binary: 011 11000
    code_group_Par[121] = 10'b1001100011; //Octect Value in Binary: 011 11001
    code_group_Par[122] = 10'b0101100011; //Octect Value in Binary: 011 11010
    code_group_Par[123] = 10'b0010011100; //Octect Value in Binary: 011 11011
    code_group_Par[124] = 10'b0011100011; //Octect Value in Binary: 011 11100
    code_group_Par[125] = 10'b0100011100; //Octect Value in Binary: 011 11101
    code_group_Par[126] = 10'b1000011100; //Octect Value in Binary: 011 11110
    code_group_Par[127] = 10'b0101001100; //Octect Value in Binary: 011 11111
    code_group_Par[128] = 10'b0110001101; //Octect Value in Binary: 100 00000
    code_group_Par[129] = 10'b1000101101; //Octect Value in Binary: 100 00001
    code_group_Par[130] = 10'b0100101101; //Octect Value in Binary: 100 00010
    code_group_Par[131] = 10'b1100010010; //Octect Value in Binary: 100 00011
    code_group_Par[132] = 10'b0010101101; //Octect Value in Binary: 100 00100
    code_group_Par[133] = 10'b1010010010; //Octect Value in Binary: 100 00101
    code_group_Par[134] = 10'b0110010010; //Octect Value in Binary: 100 00110
    code_group_Par[135] = 10'b0001110010; //Octect Value in Binary: 100 00111
    code_group_Par[136] = 10'b0001101101; //Octect Value in Binary: 100 01000
    code_group_Par[137] = 10'b1001010010; //Octect Value in Binary: 100 01001
    code_group_Par[138] = 10'b0101010010; //Octect Value in Binary: 100 01010
    code_group_Par[139] = 10'b1101000010; //Octect Value in Binary: 100 01011
    code_group_Par[140] = 10'b0011010010; //Octect Value in Binary: 100 01100
    code_group_Par[141] = 10'b1011000010; //Octect Value in Binary: 100 01101
    code_group_Par[142] = 10'b0111000010; //Octect Value in Binary: 100 01110
    code_group_Par[143] = 10'b1010001101; //Octect Value in Binary: 100 01111
    code_group_Par[144] = 10'b1001001101; //Octect Value in Binary: 100 10000
    code_group_Par[145] = 10'b1000110010; //Octect Value in Binary: 100 10001
    code_group_Par[146] = 10'b0100110010; //Octect Value in Binary: 100 10010
    code_group_Par[147] = 10'b1100100010; //Octect Value in Binary: 100 10011
    code_group_Par[148] = 10'b0010110010; //Octect Value in Binary: 100 10100
    code_group_Par[149] = 10'b1010100010; //Octect Value in Binary: 100 10101
    code_group_Par[150] = 10'b0110100010; //Octect Value in Binary: 100 10110
    code_group_Par[151] = 10'b0001011101; //Octect Value in Binary: 100 10111
    code_group_Par[152] = 10'b0011001101; //Octect Value in Binary: 100 11000
    code_group_Par[153] = 10'b1001100010; //Octect Value in Binary: 100 11001
    code_group_Par[154] = 10'b0101100010; //Octect Value in Binary: 100 11010
    code_group_Par[155] = 10'b0010011101; //Octect Value in Binary: 100 11011
    code_group_Par[156] = 10'b0011100010; //Octect Value in Binary: 100 11100
    code_group_Par[157] = 10'b0100011101; //Octect Value in Binary: 100 11101
    code_group_Par[158] = 10'b1000011101; //Octect Value in Binary: 100 11110
    code_group_Par[159] = 10'b0101001101; //Octect Value in Binary: 100 11111
    code_group_Par[160] = 10'b0110001010; //Octect Value in Binary: 101 00000
    code_group_Par[161] = 10'b1000101010; //Octect Value in Binary: 101 00001
    code_group_Par[162] = 10'b0100101010; //Octect Value in Binary: 101 00010
    code_group_Par[163] = 10'b1100011010; //Octect Value in Binary: 101 00011
    code_group_Par[164] = 10'b0010101010; //Octect Value in Binary: 101 00100
    code_group_Par[165] = 10'b1010011010; //Octect Value in Binary: 101 00101
    code_group_Par[166] = 10'b0110011010; //Octect Value in Binary: 101 00110
    code_group_Par[167] = 10'b0001111010; //Octect Value in Binary: 101 00111
    code_group_Par[168] = 10'b0001101010; //Octect Value in Binary: 101 01000
    code_group_Par[169] = 10'b1001011010; //Octect Value in Binary: 101 01001
    code_group_Par[170] = 10'b0101011010; //Octect Value in Binary: 101 01010
    code_group_Par[171] = 10'b1101001010; //Octect Value in Binary: 101 01011
    code_group_Par[172] = 10'b0011011010; //Octect Value in Binary: 101 01100
    code_group_Par[173] = 10'b1011001010; //Octect Value in Binary: 101 01101
    code_group_Par[174] = 10'b0111001010; //Octect Value in Binary: 101 01110
    code_group_Par[175] = 10'b1010001010; //Octect Value in Binary: 101 01111
    code_group_Par[176] = 10'b1001001010; //Octect Value in Binary: 101 10000
    code_group_Par[177] = 10'b1000111010; //Octect Value in Binary: 101 10001
    code_group_Par[178] = 10'b0100111010; //Octect Value in Binary: 101 10010
    code_group_Par[179] = 10'b1100101010; //Octect Value in Binary: 101 10011
    code_group_Par[180] = 10'b0010111010; //Octect Value in Binary: 101 10100
    code_group_Par[181] = 10'b1010101010; //Octect Value in Binary: 101 10101
    code_group_Par[182] = 10'b0110101010; //Octect Value in Binary: 101 10110
    code_group_Par[183] = 10'b0001011010; //Octect Value in Binary: 101 10111
    code_group_Par[184] = 10'b0011001010; //Octect Value in Binary: 101 11000
    code_group_Par[185] = 10'b1001101010; //Octect Value in Binary: 101 11001
    code_group_Par[186] = 10'b0101101010; //Octect Value in Binary: 101 11010
    code_group_Par[187] = 10'b0010011010; //Octect Value in Binary: 101 11011
    code_group_Par[188] = 10'b0011101010; //Octect Value in Binary: 101 11100
    code_group_Par[189] = 10'b0100011010; //Octect Value in Binary: 101 11101
    code_group_Par[190] = 10'b1000011010; //Octect Value in Binary: 101 11110
    code_group_Par[191] = 10'b0101001010; //Octect Value in Binary: 101 11111
    code_group_Par[192] = 10'b0110000110; //Octect Value in Binary: 110 00000
    code_group_Par[193] = 10'b1000100110; //Octect Value in Binary: 110 00001
    code_group_Par[194] = 10'b0100100110; //Octect Value in Binary: 110 00010
    code_group_Par[195] = 10'b1100010110; //Octect Value in Binary: 110 00011
    code_group_Par[196] = 10'b0010100110; //Octect Value in Binary: 110 00100
    code_group_Par[197] = 10'b1010010110; //Octect Value in Binary: 110 00101
    code_group_Par[198] = 10'b0110010110; //Octect Value in Binary: 110 00110
    code_group_Par[199] = 10'b0001110110; //Octect Value in Binary: 110 00111
    code_group_Par[200] = 10'b0001100110; //Octect Value in Binary: 110 01000
    code_group_Par[201] = 10'b1001010110; //Octect Value in Binary: 110 01001
    code_group_Par[202] = 10'b0101010110; //Octect Value in Binary: 110 01010
    code_group_Par[203] = 10'b1101000110; //Octect Value in Binary: 110 01011
    code_group_Par[204] = 10'b0011010110; //Octect Value in Binary: 110 01100
    code_group_Par[205] = 10'b1011000110; //Octect Value in Binary: 110 01101
    code_group_Par[206] = 10'b0111000110; //Octect Value in Binary: 110 01110
    code_group_Par[207] = 10'b1010000110; //Octect Value in Binary: 110 01111
    code_group_Par[208] = 10'b1001000110; //Octect Value in Binary: 110 10000
    code_group_Par[209] = 10'b1000110110; //Octect Value in Binary: 110 10001
    code_group_Par[210] = 10'b0100110110; //Octect Value in Binary: 110 10010
    code_group_Par[211] = 10'b1100100110; //Octect Value in Binary: 110 10011
    code_group_Par[212] = 10'b0010110110; //Octect Value in Binary: 110 10100
    code_group_Par[213] = 10'b1010100110; //Octect Value in Binary: 110 10101
    code_group_Par[214] = 10'b0110100110; //Octect Value in Binary: 110 10110
    code_group_Par[215] = 10'b0001010110; //Octect Value in Binary: 110 10111
    code_group_Par[216] = 10'b0011000110; //Octect Value in Binary: 110 11000
    code_group_Par[217] = 10'b1001100110; //Octect Value in Binary: 110 11001
    code_group_Par[218] = 10'b0101100110; //Octect Value in Binary: 110 11010
    code_group_Par[219] = 10'b0010010110; //Octect Value in Binary: 110 11011
    code_group_Par[220] = 10'b0011100110; //Octect Value in Binary: 110 11100
    code_group_Par[221] = 10'b0100010110; //Octect Value in Binary: 110 11101
    code_group_Par[222] = 10'b1000010110; //Octect Value in Binary: 110 11110
    code_group_Par[223] = 10'b0101000110; //Octect Value in Binary: 110 11111
    code_group_Par[224] = 10'b0110001110; //Octect Value in Binary: 111 00000
    code_group_Par[225] = 10'b1000101110; //Octect Value in Binary: 111 00001
    code_group_Par[226] = 10'b0100101110; //Octect Value in Binary: 111 00010
    code_group_Par[227] = 10'b1100010001; //Octect Value in Binary: 111 00011
    code_group_Par[228] = 10'b0010101110; //Octect Value in Binary: 111 00100
    code_group_Par[229] = 10'b1010010001; //Octect Value in Binary: 111 00101
    code_group_Par[230] = 10'b0110010001; //Octect Value in Binary: 111 00110
    code_group_Par[231] = 10'b0001110001; //Octect Value in Binary: 111 00111
    code_group_Par[232] = 10'b0001101110; //Octect Value in Binary: 111 01000
    code_group_Par[233] = 10'b1001010001; //Octect Value in Binary: 111 01001
    code_group_Par[234] = 10'b0101010001; //Octect Value in Binary: 111 01010
    code_group_Par[235] = 10'b1101001000; //Octect Value in Binary: 111 01011
    code_group_Par[236] = 10'b0011010001; //Octect Value in Binary: 111 01100
    code_group_Par[237] = 10'b1011001000; //Octect Value in Binary: 111 01101
    code_group_Par[238] = 10'b0111001000; //Octect Value in Binary: 111 01110
    code_group_Par[239] = 10'b1010001110; //Octect Value in Binary: 111 01111
    code_group_Par[240] = 10'b1001001110; //Octect Value in Binary: 111 10000
    code_group_Par[241] = 10'b1000110001; //Octect Value in Binary: 111 10001
    code_group_Par[242] = 10'b0100110001; //Octect Value in Binary: 111 10010
    code_group_Par[243] = 10'b1100100001; //Octect Value in Binary: 111 10011
    code_group_Par[244] = 10'b0010110001; //Octect Value in Binary: 111 10100
    code_group_Par[245] = 10'b1010100001; //Octect Value in Binary: 111 10101
    code_group_Par[246] = 10'b0110100001; //Octect Value in Binary: 111 10110
    code_group_Par[247] = 10'b0001011110; //Octect Value in Binary: 111 10111
    code_group_Par[248] = 10'b0011001110; //Octect Value in Binary: 111 11000
    code_group_Par[249] = 10'b1001100001; //Octect Value in Binary: 111 11001
    code_group_Par[250] = 10'b0101100001; //Octect Value in Binary: 111 11010
    code_group_Par[251] = 10'b0010011110; //Octect Value in Binary: 111 11011
    code_group_Par[252] = 10'b0011100001; //Octect Value in Binary: 111 11100
    code_group_Par[253] = 10'b0100011110; //Octect Value in Binary: 111 11101
    code_group_Par[254] = 10'b1000011110; //Octect Value in Binary: 111 11110
    code_group_Par[255] = 10'b0101001110; //Octect Value in Binary: 111 11111
    code_group_Par[256] = 10'b1100001011; //Octect Value in Binary: 000 11100
    code_group_Par[257] = 10'b1100000110; //Octect Value in Binary: 001 11100
    code_group_Par[258] = 10'b1100001010; //Octect Value in Binary: 010 11100
    code_group_Par[259] = 10'b1100001100; //Octect Value in Binary: 011 11100
    code_group_Par[260] = 10'b1100001101; //Octect Value in Binary: 100 11100
    code_group_Par[261] = 10'b1100000101; //Octect Value in Binary: 101 11100
    code_group_Par[262] = 10'b1100001001; //Octect Value in Binary: 110 11100
    code_group_Par[263] = 10'b1100000111; //Octect Value in Binary: 111 11100
    code_group_Par[264] = 10'b0001010111; //Octect Value in Binary: 111 10111
    code_group_Par[265] = 10'b0010010111; //Octect Value in Binary: 111 11011
    code_group_Par[266] = 10'b0100010111; //Octect Value in Binary: 111 11101
    code_group_Par[267] = 10'b1000010111; //Octect Value in Binary: 111 11110
    
    end
    
    
    
    
endmodule
